* Include Directives
.include '90nm_bulk.pm' MOS

* Component Definitions
M1 CLK_NOT CLK V1 V1 PMOS W=120n L=90n
M2 CLK_NOT CLK 0 0 NMOS W=150n L=90n

M3 D_NOT D V1 V1 PMOS W=120n L=90n
M4 D_NOT D 0 0 NMOS W=150n L=90n

* MASTER-SLAVE FLIP FLOP

M5 D_NOT CLK 01 V2 PMOS W=120n L=90n
M6 D_NOT CLK_NOT 01 0 NMOS W=150n L=90n

M7 D_NOT CLK 01 V2 PMOS W=120n L=90n
M8 D_NOT CLK_NOT 01 0 NMOS W=150n L=90n

M3 Y X V2 V2 PMOS W=120n L=90n
M4 Y X 0 0 NMOS W=150n L=90n
M5 OUT Y V3 V3 PMOS W=120n L=90n
M6 OUT Y 0 0 NMOS W=150n L=90n


VDD1 V1 0 1.2V
VDD2 V2 0 1.2V
VDD3 V3 0 1.2V
VDD4 V4 0 1.2V

Vd D 0 PULSE(0 2.5 0 0.1ns 0.1ns 1ns 2.2ns)
Vckl CLK 0 PULSE(0 2.5 0 0.1ns 0.1ns 1ns 2.2ns)

C1 OUT 0 0.5fF

* NG-Spice Simulation Commands
.OPTIONS NOPAGE NUMDGT=6 UNITS=Degress WIDTH=104
.PRINT TRAN V(OUT,0) V(OUT)
.TRAN 1.00n 10.00n 0.00n

.END

